
module clktrial2 (
	clk);	

	output		clk;
endmodule
