module addrpc(in1,res);
input [7:0] in1;
output [7:0] res;
assign res=in1+1;
endmodule