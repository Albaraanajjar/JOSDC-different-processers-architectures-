// clktrial2.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module clktrial2 (
		output wire  clk  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (1),
		.CLOCK_UNIT (1000)
	) clock_source_0 (
		.clk (clk)  // clk.clk
	);

endmodule
