
module clktrial1 (
	clk);	

	output		clk;
endmodule
